module Decoder32_5(
    input [4:0] decoder_in,
    output reg [31:0] decoder_out
    );
    always @(*) begin
        case (decoder_in)
        5'd0: decoder_out = 32'b00000000000000000000000000000001;
        5'd1: decoder_out = 32'b00000000000000000000000000000010;
        5'd2: decoder_out = 32'b00000000000000000000000000000100;
        5'd3: decoder_out = 32'b00000000000000000000000000001000;
        5'd4: decoder_out = 32'b00000000000000000000000000010000;
        5'd5: decoder_out = 32'b00000000000000000000000000100000;
        5'd6: decoder_out = 32'b00000000000000000000000001000000;
        5'd7: decoder_out = 32'b00000000000000000000000010000000;
        5'd8: decoder_out = 32'b00000000000000000000000100000000;
        5'd9: decoder_out = 32'b00000000000000000000001000000000;
        5'd10: decoder_out = 32'b00000000000000000000010000000000;
        5'd11: decoder_out = 32'b00000000000000000000100000000000;
        5'd12: decoder_out = 32'b00000000000000000001000000000000;
        5'd13: decoder_out = 32'b00000000000000000010000000000000;
        5'd14: decoder_out = 32'b00000000000000000100000000000000;
        5'd15: decoder_out = 32'b00000000000000001000000000000000;
        5'd16: decoder_out = 32'b00000000000000010000000000000000;
        5'd17: decoder_out = 32'b00000000000000100000000000000000;
        5'd18: decoder_out = 32'b00000000000001000000000000000000;
        5'd19: decoder_out = 32'b00000000000010000000000000000000;
        5'd20: decoder_out = 32'b00000000000100000000000000000000;
        5'd21: decoder_out = 32'b00000000001000000000000000000000;
        5'd22: decoder_out = 32'b00000000010000000000000000000000;
        5'd23: decoder_out = 32'b00000000100000000000000000000000;
        5'd24: decoder_out = 32'b00000001000000000000000000000000;
        5'd25: decoder_out = 32'b00000010000000000000000000000000;
        5'd26: decoder_out = 32'b00000100000000000000000000000000;
        5'd27: decoder_out = 32'b00001000000000000000000000000000;
        5'd28: decoder_out = 32'b00010000000000000000000000000000;
        5'd29: decoder_out = 32'b00100000000000000000000000000000;
        5'd30: decoder_out = 32'b01000000000000000000000000000000;
        default: decoder_out = 32'b10000000000000000000000000000000;
         
        endcase
    end


endmodule
